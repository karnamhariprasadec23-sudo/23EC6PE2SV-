//------------------------------------------------------------------------------
//File       : dummy_dut.sv
//Author     : karnam hariprasad saisahithi( 1BM23EC315 )
//Created    : 2026-02-24
//Module     : dummy_dut
//Project    : SystemVerilog and Verification (23EC6PE2SV)
//Faculty    : Prof. Ajaykumar Devarapalli
//Description: A placeholder dummy DUT for the class-based Packet verification lab.
//------------------------------------------------------------------------------

module dummy_dut;
endmodule
