hsef
